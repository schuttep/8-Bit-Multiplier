module Block_Sprite(
                    
					 output logic [3:0] I_0 [4],
					 output logic [3:0] I_1 [4],
					 output logic [3:0] square [4],
					 
    				 output logic [3:0] J_0 [4],
       				 output logic [3:0] J_1 [4],
    				 output logic [3:0] J_2 [4],
    				 output logic [3:0] J_3 [4],
 				 
					 output logic [3:0] T_0 [4],
					 output logic [3:0] T_1 [4],
					 output logic [3:0] T_2 [4],
					 output logic [3:0] T_3 [4],
					 
					 output logic [3:0] L_0 [4],
					 output logic [3:0] L_1 [4],
					 output logic [3:0] L_2 [4],
					 output logic [3:0] L_3 [4],
					 
					 output logic [3:0] S_0 [4],
					 output logic [3:0] S_1 [4],

					 output logic [3:0] Z_0 [4],
					 output logic [3:0] Z_1 [4]

					 );
	 
	
	always_comb	
	begin
	
	// I_0
	  I_0[0] = 4'b1111;
      I_0[1] = 4'b0000;
      I_0[2] = 4'b0000;
      I_0[3] = 4'b0000;
      
      //I_1
      I_1[0] = 4'b1000;
      I_1[1] = 4'b1000;
      I_1[2] = 4'b1000;
      I_1[3] = 4'b1000;
        
    // square
      square[0] = 4'b1100;
      square[1] = 4'b1100;
      square[2] = 4'b0000;
      square[3] = 4'b0000;
	
         
      // T_0
	  T_0[0] = 4'b0100;
      T_0[1] = 4'b1110;
      T_0[2] = 4'b0000;
      T_0[3] = 4'b0000;
         
     // T_1
      T_1[0] = 4'b1000;
      T_1[1] = 4'b1100;
      T_1[2] = 4'b1000;
      T_1[3] = 4'b0000;

    // T_2
    
      T_2[0] = 4'b1110;
      T_2[1] = 4'b0100;
      T_2[2] = 4'b0000;
      T_2[3] = 4'b0000;
      
     // T_3

      T_3[0] = 4'b0100;
      T_3[1] = 4'b1100;
      T_3[2] = 4'b0100;
      T_3[3] = 4'b0000;
      
      // J_0
      J_0[0] = 4'b1000;
      J_0[1] = 4'b1110;
      J_0[2] = 4'b0000;
      J_0[3] = 4'b0000;
      
      // J_1
      J_1[0] = 4'b1100;
      J_1[1] = 4'b1000;
      J_1[2] = 4'b1000;
      J_1[3] = 4'b0000;  
             
      // J_2
      J_2[0] = 4'b1110;
      J_2[1] = 4'b0010;
      J_2[2] = 4'b0000;
      J_2[3] = 4'b0000;       
      
      // J_3
      J_3[0] = 4'b0100;
      J_3[1] = 4'b0100;
      J_3[2] = 4'b1100;
      J_3[3] = 4'b0000;       
                                              
     // L_0
      L_0[0] = 4'b0010;
      L_0[1] = 4'b1110;
      L_0[2] = 4'b0000;
      L_0[3] = 4'b0000;
      
      // L_1
      L_1[0] = 4'b1000;
      L_1[1] = 4'b1000;
      L_1[2] = 4'b1100;
      L_1[3] = 4'b0000;  
             
      // L_2
      L_2[0] = 4'b1110;
      L_2[1] = 4'b1000;
      L_2[2] = 4'b0000;
      L_2[3] = 4'b0000;       
      
      // L_3
      L_3[0] = 4'b1100;
      L_3[1] = 4'b0100;
      L_3[2] = 4'b0100;
      L_3[3] = 4'b0000; 
      
      
      // S_0
      S_0[0] = 4'b0110;
      S_0[1] = 4'b1100;
      S_0[2] = 4'b0000;
      S_0[3] = 4'b0000;
      
      // S_1
      S_1[0] = 4'b1000;
      S_1[1] = 4'b1100;
      S_1[2] = 4'b0100;
      S_1[3] = 4'b0000;
      
      
      // Z_0
      Z_0[0] = 4'b1100;
      Z_0[1] = 4'b0110;
      Z_0[2] = 4'b0000;
      Z_0[3] = 4'b0000;
      
      // Z_1
      Z_1[0] = 4'b0100;
      Z_1[1] = 4'b1100;
      Z_1[2] = 4'b1000;
      Z_1[3] = 4'b0000;

 end
endmodule
